library verilog;
use verilog.vl_types.all;
entity g03_addr_vlg_vec_tst is
end g03_addr_vlg_vec_tst;
