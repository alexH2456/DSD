library verilog;
use verilog.vl_types.all;
entity g03_rules_test_vlg_vec_tst is
end g03_rules_test_vlg_vec_tst;
