library verilog;
use verilog.vl_types.all;
entity g02_lab5_rules_dealer_vlg_vec_tst is
end g02_lab5_rules_dealer_vlg_vec_tst;
