library verilog;
use verilog.vl_types.all;
entity g03_stack52_vlg_vec_tst is
end g03_stack52_vlg_vec_tst;
