library verilog;
use verilog.vl_types.all;
entity g03_addr_vlg_check_tst is
    port(
        Cout            : in     vl_logic;
        S0              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end g03_addr_vlg_check_tst;
