library verilog;
use verilog.vl_types.all;
entity g03_lab3_vlg_vec_tst is
end g03_lab3_vlg_vec_tst;
