library verilog;
use verilog.vl_types.all;
entity g03_lab4_vlg_check_tst is
    port(
        legal           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end g03_lab4_vlg_check_tst;
